`define     VCS_SIMULATION
