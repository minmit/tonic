`define SEND_DD_CONTEXT             1'b0
`define USER_CONTEXT_W              (3 * `FLOW_SEQ_NUM_W + `FLOW_WIN_IND_W + `FLAG_W)

`define RTO_LOW_THRESH              3
`define RTO_LOW                     500
`define RTO_HIGH                    2000


