`define   USER_CONTEXT_W          40
