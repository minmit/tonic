`define   SEND_DD_CONTEXT     1'b0
`define   USER_CONTEXT_W    (2 * `FLAG_W + 3 * `FLOW_SEQ_NUM_W + 6 * `FLOW_WIN_SIZE_W) 

`define   DUP_ACKS_THRESH               3 



