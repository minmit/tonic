`define SEND_DD_CONTEXT     1'b0
`define USER_CONTEXT_W      1
